Question 9

Vdd 1 0 10
vd 1 2 0
rd 2 3 4k
vd1 1 5 0

r1 5 4 7.5k
r2 4 0 3.2k
c1 4 6 2.2u
c2 3 8 2.2u
rl 8 0 100k
rg 6 7 1k

vin 7 0 sin (0 100m 1k 0 0 0)

M1 3 4 0 0 MN4007

.model MN4007 NMOS(Kp=500u Vto=1.5 Lambda=0.01 Gamma=0.6 Tox=1200n Phi=.6 Rs=0 Rd=0 Cbd=2.0p Cbs=2.0p Pb=.8 Cgso=0.1p Cgdo=0.1p Is=16.64p)
.tran 0.01ms 10ms 0.1ms
.control
op
run

plot v(7) v(8)
.endc
.end
