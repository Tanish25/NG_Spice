Question-2

Vcc 3 0 5V
Vgs 4 0 5V
Vd 3 1 0                                                                                                                                                                            
R1 1 2 100
M1 2 4 0 0 MN4007

.model MN4007 NMOS(Kp=500u Vto=1.5 Lambda=0.01 Gamma=0.6 Tox=1200n Phi=.6 Rs=0 Rd=0 Cbd=2.0p Cbs=2.0p Pb=.8 Cgso=0.1p Cgdo=0.1p Is=16.64p)

.dc Vcc 0.1 5 0.2 Vgs 0 5 0.2
*.tran 0.001ms 1ms
.control
run

plot i(Vd) vs v(2)
plot v(2)/i(Vd)

.endc
.end

