Common Emitter Amplifier

Vcc 3 0 12
Vin 4 0 1
Vdc 1 2 0
Vdb 5 8 0
Vde 6 9 0

.MODEL Q2N2222A NPN(IS=8.11E-14 BF=205 VAF=113 IKF=0.5 ISE=1.06E-11+ NE=2 BR=4 VAR=24 IKR=0.225 RB=1.37 RE=0.343 RC=0.137 CJE=2.95E-11+ TF=3.97E-10 CJC=1.52E-11 TR=8.5E-8 XTB=1.5)

Q1 2 8 6 Q2N2222A

Rc 3 1 5k
R1 3 5 33k
R2 5 0 10k
Re 9 0 2k

*Control Statements
.control
op
dc vin 0.01 1 0.02
run

*Plotting the output
plot i(Vdb)
plot i(Vdc)
plot i(Vde)
plot v(6)
plot v(1)


.endc
.end
