Q5
.include ua741.txt
Vin 2 3 dc 0 ac 1
R1 3 4 5k
C1 4 0 0.1u
X1 4 5 5 9 10 UA741
Vp1 9 0 dc +15V
Vm1 15 0 dc -15V
R2 5 6 5500
R3 6 7 5500
X1 0 6 UA741
R4 6 8 5500
X2 8 1 8 11 12 UA741
Vp2 11 0 dc +15V
Vm2 12 0 dc -15V
X3 6 13 14 15 7 UA741
Vp3 14 0 dc +15V
vm3 15 0 dc -15V 
.tran 0.001ms 1ms uic
.control
run
plot ac v(7)
.endc
.end